-- This file is part of easyFPGA.
-- Copyright 2013,2014 os-cillation GmbH
--
-- easyFPGA is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- easyFPGA is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with easyFPGA.  If not, see <http://www.gnu.org/licenses/>.

-------------------------------------------------------------------------------
-- P A R T    N A M E
-- (<name>.vhd)
--
-- Structural
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

-------------------------------------------------------------------------------
ENTITY <name> is
-------------------------------------------------------------------------------
   port (
   );
end <name>;

-------------------------------------------------------------------------------
ARCHITECTURE structural of <name> is
-------------------------------------------------------------------------------
   ----------------------------------------------
   -- constants
   ----------------------------------------------

   ----------------------------------------------
   -- signals
   ----------------------------------------------

--------------------------------------------------------------------------------
begin -- architecture structural
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
INSTANCE_A : entity work.test234
-------------------------------------------------------------------------------
   port map (
   );

end structural;
